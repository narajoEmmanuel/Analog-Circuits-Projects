Proyecto_Laboratorio_Electronica_Potencia
 *Ciclo convertidor Trif�sico - Monof�sico
 *Estudiantes:
 		*Jose Fabio Navarro Naranjo 2019049626
 		*Emmanuel Naranjo Blanco   2019053605
 		*Adrian Dittel Retana             2019007945
 
*Definicion de parametros para la simulacion del circuito

*Entradas
.param V_in={120};  *Tension RMS de entrada por fase
.param f_in={260} ; *Frecuencia de entrada (entre 120Hz y 400Hz)
.param f_out={65} ;*Frecuencia de salida (entre 30Hz y 100Hz))
.param alfa={131}; *Angulo de disparo
.param carga={82.3} ;*carga a alimentar (resistiva)

*Derivaciones de las entradas
.param V_pico={V_in*sqrt(2)}; *Tension pico en la entrada
.param delay_p={alfa/(360*f_in)}; *Delay para la fase P
.param delay_n={(periodo_in/2)+delay_p}; *Delay para la fase N
.param pw={1/(3*f_in)}; *Tiempo en alto de los SCR (pulse width) 
.param periodo_in={1/f_in}; *Periodo de la se�al de entrada
.param periodo_out={1/f_out}; *Periodo de la se�al de salida
.param pw_pn={0.5*periodo_out}; *Tiempo en alto de las se�ales p y n

*Componentes del circuito

*Definicion de las entradas de fase 
Van 1 0 Sin(0 {V_pico} {f_in} 0 0 -30); *fase A
Vbn 2 0 Sin(0 {V_pico} {f_in} 0 0 -150); *fase B
Vcn 3 0 Sin(0 {V_pico} {f_in} 0 0 -270); *fase C

*Para la implemetacion de los SCR se van a utilizar diodos en combinacion con switches que en conjunto simulan el comportamiento deseado

*P Converter (Switches y Diodos)

sw1p 1 4 18 0 smod
dio1p 4 5 dmod

sw3p 2 6 19 0 smod
dio3p 6 5 dmod

sw5p 3 7 20 0 smod
dio5p 7 5 dmod

sw2p 8 9 21 0 smod
dio2p 9 1 dmod

sw4p 8 10 22 0 smod
dio4p 10 2 dmod

sw6p 8 11 23 0 smod
dio6p 11 3 dmod

*N Converter (Switches y Diodos)

sw1n 5 12 24 0 smod
dio1n 12 1 dmod

sw3n 5 13 25 0 smod
dio3n 13 2 dmod

sw5n 5 14 26 0  smod
dio5n 14 3 dmod

sw2n 1 15 27 0 smod
dio2n 15 8 dmod

sw4n 2 16 28 0 smod
dio4n 16 8 dmod

sw6n 3 17 29 0 smod
dio6n 17 8 dmod

*Carga
r_load 5 8 {carga} 

*Control para los switches

*Control P

v1p 18 30 pulse(-5 5 {delay_p} 1ns 1ns {pw} {periodo_in})
v3p 19 30 pulse(-5 5 {delay_p + periodo_in/3} 1ns 1ns {pw} {periodo_in})
v5p 20 30 pulse(-5 5 {delay_p + 2*periodo_in/3} 1ns 1ns {pw} {periodo_in})
v2p 21 30 pulse(-5 5 {delay_p + periodo_in/2} 1ns 1ns {pw} {periodo_in})
v4p 22 30 pulse(-5 5 {delay_p + 5*periodo_in/6} 1ns 1ns {pw} {periodo_in})
v6p 23 30 pulse(-5 5 {delay_p + periodo_in/6} 1ns 1ns {pw} {periodo_in})

vc_p 30 0 pulse(5 -5 0 1ns 1ns {pw_pn} {periodo_out}); *fuente para controlar la fase P

*Control N

v1n 24 31 pulse(-5 5 {delay_n} 1ns 1ns {pw} {periodo_in})
v3n 25 31 pulse(-5 5 {delay_n + periodo_in/3} 1ns 1ns {pw} {periodo_in})
v5n 26 31 pulse(-5 5 {delay_n + 2*periodo_in/3} 1ns 1ns {pw} {periodo_in})
v2n 27 31 pulse(-5 5 {delay_n + periodo_in/2} 1ns 1ns {pw} {periodo_in})
v4n 28 31 pulse(-5 5 {delay_n + 5*periodo_in/6} 1ns 1ns {pw} {periodo_in})
v6n 29 31 pulse(-5 5 {delay_n + periodo_in/6} 1ns 1ns {pw} {periodo_in})

vc_n 31 0 pulse(5 -5 {periodo_out/2} 1ns 1ns {pw_pn} {periodo_out}); *fuente para controlar la fase N

.model smod VSWITCH(Ron=0.001m)
.model dmod d
.tran .1ms 400ms 0ms .1ms uic
*.FOUR {f_out} 30 V(5,8)
.FOUR {f_in} 30 I(Van)
.probe
.end